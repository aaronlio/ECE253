module part3(Clock, Reset, Go, Divisor, Dividend, Quotient, Remainder, ResultValid);
